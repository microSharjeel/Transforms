module HEVC_DCT32_ROM (
input  logic [4:0] row,
input  logic [4:0] col,
output logic signed [7:0] coeff
);
logic signed [7:0] COEFFS [0:31][0:31] = '{
'{ 64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64,  64},
'{ 90,  90,  90,  90,  89,  88,  87,  85,  83,  82,  80,  78,  75,  73,  70,  67,  64,  61,  57,  54,  50,  46,  43,  38,  36,  31,  25,  22,  18,  13,   9,   4},
'{ 90,  90,  90,  90,  87,  80,  70,  57,  43,  25,   9,  -9, -25, -43, -57, -70, -80, -87, -90, -90, -90, -90, -87, -80, -70, -57, -43, -25,  -9,   9,  25,  43},
'{ 90,  90,  88,  85,  82,  78,  73,  67,  61,  54,  46,  38,  31,  22,  13,   4,  -4, -13, -22, -31, -38, -46, -54, -61, -67, -73, -78, -82, -85, -88, -90, -90},
'{ 90,  90,  90,  90,  83,  67,  46,  22,  -4, -31, -54, -73, -85, -90, -88, -78, -61, -38, -13,  13,  38,  61,  78,  88,  90,  85,  73,  54,  31,   4, -22, -46},
'{ 90,  90,  87,  82,  75,  67,  57,  46,  36,  22,   9,  -4, -18, -31, -43, -54, -64, -73, -80, -85, -89, -90, -90, -88, -85, -80, -73, -64, -54, -43, -31, -18},
'{ 90,  89,  87,  83,  78,  70,  61,  50,  38,  25,  13,   0, -13, -25, -38, -50, -61, -70, -78, -83, -87, -89, -90, -89, -87, -83, -78, -70, -61, -50, -38, -25},
'{ 90,  88,  85,  78,  70,  57,  43,  25,   9,  -9, -25, -43, -57, -70, -78, -85, -88, -90, -88, -85, -78, -70, -57, -43, -25,  -9,   9,  25,  43,  57,  70,  78},
'{ 90,  90,  90,  90,  78,  54,  22, -13, -46, -73, -90, -90, -78, -54, -22,  13,  46,  73,  90,  90,  78,  54,  22, -13, -46, -73, -90, -90, -78, -54, -22,  13},
'{ 90,  88,  82,  73,  61,  46,  31,  13,  -4, -22, -38, -54, -67, -78, -85, -90, -90, -88, -82, -73, -61, -46, -31, -13,   4,  22,  38,  54,  67,  78,  85,  90},
'{ 90,  87,  80,  67,  50,  31,   9, -13, -36, -54, -70, -82, -90, -90, -85, -75, -61, -43, -22,   0,  22,  43,  61,  75,  85,  90,  90,  82,  70,  54,  36,  13},
'{ 90,  85,  73,  54,  31,   4, -22, -46, -67, -83, -90, -88, -78, -61, -38, -13,  13,  38,  61,  78,  88,  90,  83,  67,  46,  22,  -4, -31, -54, -73, -85, -90},
'{ 89,  83,  70,  50,  25,  -4, -36, -64, -85, -95, -95, -85, -64, -36,  -4,  25,  50,  70,  83,  89,  89,  83,  70,  50,  25,  -4, -36, -64, -85, -95, -95, -85},
'{ 90,  82,  67,  46,  22,  -4, -31, -54, -73, -85, -90, -88, -78, -61, -38, -13,  13,  38,  61,  78,  88,  90,  85,  73,  54,  31,   4, -22, -46, -67, -82, -90},
'{ 90,  80,  61,  36,   9, -18, -43, -64, -80, -90, -90, -80, -61, -36,  -9,  18,  43,  64,  80,  90,  90,  80,  61,  36,   9, -18, -43, -64, -80, -90, -90, -80},
'{ 90,  78,  54,  22, -13, -46, -73, -90, -90, -78, -54, -22,  13,  46,  73,  90,  90,  78,  54,  22, -13, -46, -73, -90, -90, -78, -54, -22,  13,  46,  73,  90},
'{ 89,  75,  50,  18, -18, -50, -75, -89, -89, -75, -50, -18,  18,  50,  75,  89,  89,  75,  50,  18, -18, -50, -75, -89, -89, -75, -50, -18,  18,  50,  75,  89},
'{ 90,  73,  38,  -4, -46, -82, -90, -78, -46,  -4,  38,  73,  90,  82,  46,   4, -38, -73, -90, -82, -46,  -4,  38,  73,  90,  82,  46,   4, -38, -73, -90, -82},
'{ 90,  70,  25, -25, -70, -90, -90, -70, -25,  25,  70,  90,  90,  70,  25, -25, -70, -90, -90, -70, -25,  25,  70,  90,  90,  70,  25, -25, -70, -90, -90, -70},
'{ 90,  67,  13, -46, -85, -90, -61,  -4,  54,  88,  90,  54,  -4, -61, -90, -85, -46,  13,  67,  90,  85,  46, -13, -67, -90, -85, -46,  13,  67,  90,  85,  46},
'{ 88,  61,   4, -54, -90, -85, -31,  31,  85,  90,  54,  -4, -61, -88, -88, -61,  -4,  54,  90,  85,  31, -31, -85, -90, -54,   4,  61,  88,  88,  61,   4, -54},
'{ 87,  54,  -9, -70, -90, -70,  -9,  54,  87,  87,  54,  -9, -70, -90, -70,  -9,  54,  87,  87,  54,  -9, -70, -90, -70,  -9,  54,  87,  87,  54,  -9, -70, -90},
'{ 85,  46, -22, -82, -90, -54,  13,  73,  90,  67,   4, -61, -90, -78, -31,  38,  88,  90,  54, -18, -80, -90, -50,  25,  83,  90,  46, -36, -87, -83, -22,  57},
'{ 83,  36, -36, -83, -83, -36,  36,  83,  83,  36, -36, -83, -83, -36,  36,  83,  83,  36, -36, -83, -83, -36,  36,  83,  83,  36, -36, -83, -83, -36,  36,  83},
'{ 82,  22, -54, -90, -61,  13,  78,  85,  31, -46, -90, -67,   4,  73,  88,  38, -38, -88, -73,  -4,  67,  90,  46, -31, -85, -78, -13,  61,  90,  54, -22, -82},
'{ 80,   9, -70, -87, -25,  57,  90,  43, -43, -90, -57,  25,  87,  70,  -9, -80, -80,  -9,  70,  87,  25, -57, -90, -43,  43,  90,  57, -25, -87, -70,   9,  80},
'{ 78,  -4, -82, -73,  13,  85,  67, -22, -88, -61,  31,  90,  54, -38, -90, -46,  46,  90,  38, -54, -90, -31,  61,  88,  22, -67, -85, -13,  73,  82,   4, -78},
'{ 75, -18, -89, -50,  50,  89,  18, -75, -75,  18,  89,  50, -50, -89, -18,  75,  75, -18, -89, -50,  50,  89,  18, -75, -75,  18,  89,  50, -50, -89, -18,  75},
'{ 73, -31, -90, -22,  78,  67, -38, -90, -13,  82,  61, -46, -88,  -4,  85,  54, -54, -85,   4,  88,  46, -61, -82,  13,  90,  38, -67, -78,  22,  90,  31, -73},
'{ 70, -43, -87,   9,  90,  25, -80, -57,  57,  80, -25, -90,  -9,  87,  43, -70, -70,  43,  87,  -9, -90, -25,  80,  57, -57, -80,  25,  90,   9, -87, -43,  70},
'{ 67, -54, -78,  38,  85, -22, -90,   4,  90,  13, -88, -31,  82,  46, -73, -61,  61,  73, -46, -82,  31,  88, -13, -90,  -4,  90,  22, -85, -38,  78,  54, -67},
'{ 64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64,  64, -64, -64,  64}
};
assign coeff = COEFFS[row][col];
endmodule