module HEVC_DCT8_ROM (
input  logic [2:0] row,
input  logic [2:0] col,
output logic signed [7:0] coeff  
);
logic signed [7:0] COEFFS [0:7][0:7] = '{
'{ 64,  64,  64,  64,  64,  64,  64,  64},
'{ 89,  75,  50,  18, -18, -50, -75, -89},
'{ 83,  36, -36, -83, -83, -36,  36,  83},
'{ 75, -18, -89, -50,  50,  89,  18, -75},
'{ 64, -64, -64,  64,  64, -64, -64,  64},
'{ 50, -89,  18,  75, -75, -18,  89, -50},
'{ 36, -83,  83, -36, -36,  83, -83,  36},
'{ 18, -50,  75, -89,  89, -75,  50, -18}
};
assign coeff = COEFFS[row][col];
endmodule